`include "idli_pkg.svh"


// Top-level module for the core. This is what is instantiated in the bench
// and what should eventually be used as the module in Tiny Tapeout.
module idli_top_m import idli_pkg::*; (
  // Clock and reset.
  input  var logic      i_top_gck,
  input  var logic      i_top_rst_n,

  // Low memory interface.
  output var logic      o_top_mem_lo_sck,
  output var logic      o_top_mem_lo_cs,
  input  var slice_t    i_top_mem_lo_sio,
  output var slice_t    o_top_mem_lo_sio,
  output var logic      o_top_mem_lo_en,

  // High memory interface.
  output var logic      o_top_mem_hi_sck,
  output var logic      o_top_mem_hi_cs,
  input  var slice_t    i_top_mem_hi_sio,
  output var slice_t    o_top_mem_hi_sio,
  output var logic      o_top_mem_hi_en,

  // UART interface.
  input  var logic      i_top_uart_rx,
  output var logic      o_top_uart_tx,

  // Input and output pin interface.
  input  var io_pins_t  i_top_io_pins,
  output var io_pins_t  o_top_io_pins,

  // Debug probes for the bench.
  output var debug_t    o_top_debug
);

  data_t  instr;
  logic   instr_vld;
  slice_t mem_data;
  logic   ex_redirect;
  slice_t ex_data;
  logic   ex_stall;
  logic   ex_mem_wr;
  logic   wr_acp;

  slice_t utx_data;
  logic   utx_vld;
  logic   utx_acp;

  slice_t urx_data;
  logic   urx_vld;
  logic   urx_acp;

  // TODO Move the counter into the sync/control block.
  ctr_t ctr_q;
  always_ff @(posedge i_top_gck, negedge i_top_rst_n) begin
    if (!i_top_rst_n) ctr_q <= '0;
    else              ctr_q <= ctr_q + 2'b1;
  end

always_comb o_top_debug.ctr = ctr_q;


  idli_sqi_m sqi_u (
    .i_sqi_gck        (i_top_gck),
    .i_sqi_rst_n      (i_top_rst_n),

    .i_sqi_ctr        (ctr_q),
    .i_sqi_redirect   (ex_redirect),
    .i_sqi_wr_en      (ex_mem_wr),
    .i_sqi_stall      (ex_stall),

    .i_sqi_slice      (ex_data),
    .o_sqi_slice      (mem_data),
    .o_sqi_instr      (instr),
    .o_sqi_instr_vld  (instr_vld),
    .o_sqi_wr_acp     (wr_acp),

    .o_sqi_lo_sck     (o_top_mem_lo_sck),
    .o_sqi_lo_cs      (o_top_mem_lo_cs),
    .i_sqi_lo_sio     (i_top_mem_lo_sio),
    .o_sqi_lo_sio     (o_top_mem_lo_sio),
    .o_sqi_lo_en      (o_top_mem_lo_en),

    .o_sqi_hi_sck     (o_top_mem_hi_sck),
    .o_sqi_hi_cs      (o_top_mem_hi_cs),
    .i_sqi_hi_sio     (i_top_mem_hi_sio),
    .o_sqi_hi_sio     (o_top_mem_hi_sio),
    .o_sqi_hi_en      (o_top_mem_hi_en)
  );


  idli_ex_m ex_u (
    .i_ex_gck       (i_top_gck),
    .i_ex_rst_n     (i_top_rst_n),

    .i_ex_ctr       (ctr_q),
    .i_ex_enc       (instr),
    .i_ex_enc_vld   (instr_vld),
    .i_ex_data      (mem_data),

    .o_ex_redirect  (ex_redirect),
    .o_ex_data      (ex_data),
    .o_ex_stall     (ex_stall),
    .o_ex_mem_wr    (ex_mem_wr),
    .i_ex_mem_acp   (wr_acp),

    .o_ex_utx_data  (utx_data),
    .o_ex_utx_vld   (utx_vld),
    .i_ex_utx_acp   (utx_acp),

    .i_ex_urx_data  (urx_data),
    .i_ex_urx_vld   (urx_vld),
    .o_ex_urx_acp   (urx_acp),

    .i_ex_io_pins   (i_top_io_pins),
    .o_ex_io_pins   (o_top_io_pins),

    .o_ex_debug     (o_top_debug.ex)
  );


  idli_utx_m utx_u (
    .i_utx_gck    (i_top_gck),
    .i_utx_rst_n  (i_top_rst_n),

    .i_utx_ctr    (ctr_q),
    .i_utx_data   (utx_data),
    .i_utx_vld    (utx_vld),
    .o_utx_acp    (utx_acp),

    .o_utx_data   (o_top_uart_tx)
  );


  idli_urx_m urx_u (
    .i_urx_gck    (i_top_gck),
    .i_urx_rst_n  (i_top_rst_n),

    .i_urx_ctr    (ctr_q),
    .o_urx_data   (urx_data),
    .o_urx_vld    (urx_vld),
    .i_urx_acp    (urx_acp),

    .i_urx_data   (i_top_uart_rx),

    .o_urx_debug  (o_top_debug.urx)
  );

endmodule
