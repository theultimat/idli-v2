// Wrapper for the top module for debug.
module idli_tb_m();

  // Clock and reset signals.
  logic gck;
  logic rst_n;

endmodule
